module zeroExtend (
    input logic [3:0] label,
    output logic [15:0] ZeroExtLabel
);
    assign ZeroExtLabel = { 12'b0, label };
endmodule

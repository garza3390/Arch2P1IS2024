module sbox_rom_comb (
    input  logic [7:0] address,   // Dirección de entrada (byte a sustituir)
    output logic [7:0] q          // Salida (byte sustituido)
);

    // ROM combinacional utilizando un bloque always_comb
    always_comb begin
        case (address)
            8'h00: q = 8'h63;
            8'h01: q = 8'h7C;
            8'h02: q = 8'h77;
            8'h03: q = 8'h7B;
            8'h04: q = 8'hF2;
            8'h05: q = 8'h6B;
            8'h06: q = 8'h6F;
            8'h07: q = 8'hC5;
            8'h08: q = 8'h30;
            8'h09: q = 8'h01;
            8'h0A: q = 8'h67;
            8'h0B: q = 8'h2B;
            8'h0C: q = 8'hFE;
            8'h0D: q = 8'hD7;
            8'h0E: q = 8'hAB;
            8'h0F: q = 8'h76;
            8'h10: q = 8'hCA;
            8'h11: q = 8'h82;
            8'h12: q = 8'hC9;
            8'h13: q = 8'h7D;
            8'h14: q = 8'hFA;
            8'h15: q = 8'h59;
            8'h16: q = 8'h47;
            8'h17: q = 8'hF0;
            8'h18: q = 8'hAD;
            8'h19: q = 8'hD4;
            8'h1A: q = 8'hA2;
            8'h1B: q = 8'hAF;
            8'h1C: q = 8'h9C;
            8'h1D: q = 8'hA4;
            8'h1E: q = 8'h72;
            8'h1F: q = 8'hC0;
            8'h20: q = 8'hB7;
            8'h21: q = 8'hFD;
            8'h22: q = 8'h93;
            8'h23: q = 8'h26;
            8'h24: q = 8'h36;
            8'h25: q = 8'h3F;
            8'h26: q = 8'hF7;
            8'h27: q = 8'hCC;
            8'h28: q = 8'h34;
            8'h29: q = 8'hA5;
            8'h2A: q = 8'hE5;
            8'h2B: q = 8'hF1;
            8'h2C: q = 8'h71;
            8'h2D: q = 8'hD8;
            8'h2E: q = 8'h31;
            8'h2F: q = 8'h15;
            8'h30: q = 8'h04;
            8'h31: q = 8'hC7;
            8'h32: q = 8'h23;
            8'h33: q = 8'hC3;
            8'h34: q = 8'h18;
            8'h35: q = 8'h96;
            8'h36: q = 8'h05;
            8'h37: q = 8'h9A;
            8'h38: q = 8'h07;
            8'h39: q = 8'h12;
            8'h3A: q = 8'h80;
            8'h3B: q = 8'hE2;
            8'h3C: q = 8'hEB;
            8'h3D: q = 8'h27;
            8'h3E: q = 8'hB2;
            8'h3F: q = 8'h75;
            8'h40: q = 8'h09;
            8'h41: q = 8'h83;
            8'h42: q = 8'h2C;
            8'h43: q = 8'h1A;
            8'h44: q = 8'h1B;
            8'h45: q = 8'h6E;
            8'h46: q = 8'h5A;
            8'h47: q = 8'hA0;
            8'h48: q = 8'h52;
            8'h49: q = 8'h3B;
            8'h4A: q = 8'hD6;
            8'h4B: q = 8'hB3;
            8'h4C: q = 8'h29;
            8'h4D: q = 8'hE3;
            8'h4E: q = 8'h2F;
            8'h4F: q = 8'h84;
            8'h50: q = 8'h53;
            8'h51: q = 8'hD1;
            8'h52: q = 8'h00;
            8'h53: q = 8'hED;
            8'h54: q = 8'h20;
            8'h55: q = 8'hFC;
            8'h56: q = 8'hB1;
            8'h57: q = 8'h5B;
            8'h58: q = 8'h6A;
            8'h59: q = 8'hCB;
            8'h5A: q = 8'hBE;
            8'h5B: q = 8'h39;
            8'h5C: q = 8'h4A;
            8'h5D: q = 8'h4C;
            8'h5E: q = 8'h58;
            8'h5F: q = 8'hCF;
            8'h60: q = 8'hD0;
            8'h61: q = 8'hEF;
            8'h62: q = 8'hAA;
            8'h63: q = 8'hFB;
            8'h64: q = 8'h43;
            8'h65: q = 8'h4D;
            8'h66: q = 8'h33;
            8'h67: q = 8'h85;
            8'h68: q = 8'h45;
            8'h69: q = 8'hF9;
            8'h6A: q = 8'h02;
            8'h6B: q = 8'h7F;
            8'h6C: q = 8'h50;
            8'h6D: q = 8'h3C;
            8'h6E: q = 8'h9F;
            8'h6F: q = 8'hA8;
            8'h70: q = 8'h51;
            8'h71: q = 8'hA3;
            8'h72: q = 8'h40;
            8'h73: q = 8'h8F;
            8'h74: q = 8'h92;
            8'h75: q = 8'h9D;
            8'h76: q = 8'h38;
            8'h77: q = 8'hF5;
            8'h78: q = 8'hBC;
            8'h79: q = 8'hB6;
            8'h7A: q = 8'hDA;
            8'h7B: q = 8'h21;
            8'h7C: q = 8'h10;
            8'h7D: q = 8'hFF;
            8'h7E: q = 8'hF3;
            8'h7F: q = 8'hD2;
            8'h80: q = 8'hCD;
            8'h81: q = 8'h0C;
            8'h82: q = 8'h13;
            8'h83: q = 8'hEC;
            8'h84: q = 8'h5F;
            8'h85: q = 8'h97;
            8'h86: q = 8'h44;
            8'h87: q = 8'h17;
            8'h88: q = 8'hC4;
            8'h89: q = 8'hA7;
            8'h8A: q = 8'h7E;
            8'h8B: q = 8'h3D;
            8'h8C: q = 8'h64;
            8'h8D: q = 8'h5D;
            8'h8E: q = 8'h19;
            8'h8F: q = 8'h73;
            8'h90: q = 8'h60;
            8'h91: q = 8'h81;
            8'h92: q = 8'h4F;
            8'h93: q = 8'hDC;
            8'h94: q = 8'h22;
            8'h95: q = 8'h2A;
            8'h96: q = 8'h90;
            8'h97: q = 8'h88;
            8'h98: q = 8'h46;
            8'h99: q = 8'hEE;
            8'h9A: q = 8'hB8;
            8'h9B: q = 8'h14;
            8'h9C: q = 8'hDE;
            8'h9D: q = 8'h5E;
            8'h9E: q = 8'h0B;
            8'h9F: q = 8'hDB;
            8'hA0: q = 8'hE0;
            8'hA1: q = 8'h32;
            8'hA2: q = 8'h3A;
            8'hA3: q = 8'h0A;
            8'hA4: q = 8'h49;
            8'hA5: q = 8'h06;
            8'hA6: q = 8'h24;
            8'hA7: q = 8'h5C;
            8'hA8: q = 8'hC2;
            8'hA9: q = 8'hD3;
            8'hAA: q = 8'hAC;
            8'hAB: q = 8'h62;
            8'hAC: q = 8'h91;
            8'hAD: q = 8'h95;
            8'hAE: q = 8'hE4;
            8'hAF: q = 8'h79;
            8'hB0: q = 8'hE7;
            8'hB1: q = 8'hC8;
            8'hB2: q = 8'h37;
            8'hB3: q = 8'h6D;
            8'hB4: q = 8'h8D;
            8'hB5: q = 8'hD5;
            8'hB6: q = 8'h4E;
            8'hB7: q = 8'hA9;
            8'hB8: q = 8'h6C;
            8'hB9: q = 8'h56;
            8'hBA: q = 8'hF4;
            8'hBB: q = 8'hEA;
            8'hBC: q = 8'h65;
            8'hBD: q = 8'h7A;
            8'hBE: q = 8'hAE;
            8'hBF: q = 8'h08;
            8'hC0: q = 8'hBA;
            8'hC1: q = 8'h78;
            8'hC2: q = 8'h25;
            8'hC3: q = 8'h2E;
            8'hC4: q = 8'h1C;
            8'hC5: q = 8'hA6;
            8'hC6: q = 8'hB4;
            8'hC7: q = 8'hC6;
            8'hC8: q = 8'hE8;
            8'hC9: q = 8'hDD;
            8'hCA: q = 8'h74;
            8'hCB: q = 8'h1F;
            8'hCC: q = 8'h4B;
            8'hCD: q = 8'hBD;
            8'hCE: q = 8'h8B;
            8'hCF: q = 8'h8A;
            8'hD0: q = 8'h70;
            8'hD1: q = 8'h3E;
            8'hD2: q = 8'hB5;
            8'hD3: q = 8'h66;
            8'hD4: q = 8'h48;
            8'hD5: q = 8'h03;
            8'hD6: q = 8'hF6;
            8'hD7: q = 8'h0E;
            8'hD8: q = 8'h61;
            8'hD9: q = 8'h35;
            8'hDA: q = 8'h57;
            8'hDB: q = 8'hB9;
            8'hDC: q = 8'h86;
            8'hDD: q = 8'hC1;
            8'hDE: q = 8'h1D;
            8'hDF: q = 8'h9E;
            8'hE0: q = 8'hE1;
            8'hE1: q = 8'hF8;
            8'hE2: q = 8'h98;
            8'hE3: q = 8'h11;
            8'hE4: q = 8'h69;
            8'hE5: q = 8'hD9;
            8'hE6: q = 8'h8E;
            8'hE7: q = 8'h94;
            8'hE8: q = 8'h9B;
            8'hE9: q = 8'h1E;
            8'hEA: q = 8'h87;
            8'hEB: q = 8'hE9;
            8'hEC: q = 8'hCE;
            8'hED: q = 8'h55;
            8'hEE: q = 8'h28;
            8'hEF: q = 8'hDF;
            8'hF0: q = 8'h8C;
            8'hF1: q = 8'hA1;
            8'hF2: q = 8'h89;
            8'hF3: q = 8'h0D;
            8'hF4: q = 8'hBF;
            8'hF5: q = 8'hE6;
            8'hF6: q = 8'h42;
            8'hF7: q = 8'h68;
            8'hF8: q = 8'h41;
            8'hF9: q = 8'h99;
            8'hFA: q = 8'h2D;
            8'hFB: q = 8'h0F;
            8'hFC: q = 8'hB0;
            8'hFD: q = 8'h54;
            8'hFE: q = 8'hBB;
            8'hFF: q = 8'h16;
            default: q = 8'h00;
        endcase
    end

endmodule

module adder (input logic [15:0] a, b,
				  output logic [15:0] y
);

	assign y = a + b;
	
endmodule